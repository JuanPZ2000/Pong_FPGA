LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY romRed2 IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=320;
					ADDR_WIDTH	:	INTEGER:=8);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF romRed2 IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111000000000000000000111111111100111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111100000000000000000011111111111110011111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111000000000000000001111111111111111100111111111111111111111111111111111111111111111111111111111100000000011111111111111111111000001111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111110000000000000000111111111111111111110011111111111111111111111111111111111111111111111111111111111100000011111111111111111000111111111111111111110000100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111000000000000000011111111111111111111111001111111111111111111111111111111111111111111111111111111111110000011111111111111100111111111111111111111110000000111110100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111110000000000000001111111111111111111111111100111111111111111111111111111111111111111111111111111111111111000001111111111110011111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111100000000000000011111111111111111111111111110011111111111111111111111111111111111111111111111111111111111000000111111111001111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111100000000000000111111111111111111111111111111011111111111111111111111111111111111111111111111111111111110000000011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111110011100000000011111111111111111111111111111111101111111111111111111111111111111111111111111111111111111110000000011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111100001110000000111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111100000000011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111000001111000001111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111100000000011100111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111000000111100011111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111000000000011011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111110000000001110111111111111111111111000000000111111111101111111111111111111111111111111111111111111111111111100000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111110001000000011111111111111111111100000000000001111111110111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111110111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111000010000000001111111111111111100000000000000000011111110011111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111110111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111000010000000011111111111111100000000000000000000000111111011111111111111111111111111111111111111111111111111111000000011111001111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111110000001100000011111111111110000000000000000000000000011111001111111111111111111111111111111111111111111111100000000000111111011111111111111111111111111111111111111111111111111111011111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111110000000011000111111111111100000000000000000000000000001111101111111111111111111111111111111111111111111111101111000001111111011111111111111111111111111111111111111111111111111111001111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111100000000000001111111111110000000000000000000000000000000011100111111111111111111111111111111111111111111111011111110001111110111111111111111111111111111111111111111111111111111111001111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111000000000000011111111111111000000000000000000000000000000001110111111111111111111111111111111111111111111111111111111001110000111111111111111111111111101111111111111111111111111111010111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111000000000000011111111110111100000000000000000000000000000000111011111111111111111111111111111111111111111111111101111000000000111111111111111111111111001111111111111111111111111111111011100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111110000000000000011111111000001110000000000000000000000000000000011011111111111111111111111111111111111111111110111000111000000000101100000000011101111111011111111111111111111111111111101001110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111110000000000000111111110000000111100000000000000000000000000000001001111111111111111111111111111111111111111111111000010000000001101000000000011000000110011111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111110000000000001111111110000000011110000000000000000000000000000000001111111111111111111111111111111111111111111111000010000000001000000000000011000000110110011111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111100000000000001111110011100000000111000000000000000000000000000000001111111111111111111111111111111111111111101110000000000000000000000000000000000000100100000001111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111100000000000011111100001110000000011100000000000000000000000000000000111111111111111111111111111111111111111111110000000000000010000000000000000000000001000000000000111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111000000000000011111000000111000000001110000000000000000000000000000000111111111111111111111111111111111111111011110000000000000000000000000000000000000001000000000000000011111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111000000000000011110000000001110000000011100000000000000000000000000000111111111111111111111111111111111111111011110000000000000000000000000000000000000001000000000000000000111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111110000000000000111100000000000111000000001110000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000010000000000000000000001111011111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111110000000000000111000000000000011110000000111000000000000000000000000000011111111111111111111111111111111111110111100000000000000000000110000000000000000010000000000000000000000110011111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000001110000000000000000111000000001100000000000000000000000000011111111111111111111111111111111111111111100110000000000001100110000000000000000100000000000000000000000100001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000001100000000000000000011100000000110000000000000000000000000011111111111111111111111111111111111111111100110000000000011001110000000000110000100001000000000000000000000001101111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000011000000000000000000000111000000001000000000000000000000000011111111111111111111111111111111111101111001110000000000011001100000000010110000000011000000000000000000000000000001111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000010000000000000000000000011100000000000000000000000000000000011111111111111111111111111111111111101111001111000000000111001100000000111110000000010000000000000000000000000000000001100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000001111000000000000000000000000000000001111111111111111111111111111111111011111001111000110001111011100100000111111001000110000000000000000000000000000000001000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000011100000000000000000000000000000001111111111111111111111111111111111011111011111000110001111111101100000111111001000111001011000000000000010000000000001000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000001111000000000000000000000000000001111111111111111111111111111111111011110011110000010011111111111000001111111000001111111111111100000000110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000011100000000000000000000000000001111111111111111111111111111111111111110011110000110011111111111000001111110010011111111111111111000001100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000001110000000000000000000000000001111111111111111111111111111111110111110111110000100111111111111000011111110000011111111111111111000011100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000111100000000000000000000000001111111111111111111111111111111110111100111110000100111111111111000011111110000111111111111111110000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000001110000000000000000000000001111111111111111111111111111111111111100111100000001111111111111000011111100100111111111111111110001111001000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000111100000000000000000000001111111111111111111111111111111101111101111100000001111111111111000111111100101111111111111111100011111011101000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000001110000000000000000000001111111111111111111111111111111101111101111100000001111111111111000111111000001111111111111111100111110011101000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000111000000000000000000001111111111111111111111111111111111111001111100000011111111111111000111110000011111111111111111001111110111011000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000100000000000000000000000000000000000000000000000000001110000000000000000000111111111111111111111111111111011111011111000000011111111111110000111100000011111111111111110011111110111011000110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000011110000000000000000000000000000000000000000000000000111000000000000000000111111111111111111111111111111011111011111000000011111111111110001111100000011111111111111100111111100110011001110001000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000110000000000000000000000000000000000000000000000000011100000000000000000111111111111111111111111111111011111011111000000111111111111110001111101100111111111111110011111111101110111101110001100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000100000000000000000000000000000000000000000000000000111000000000000000111111111111111111111111111111111111011111000000111111111111110001111001100111111111111100111111111001101111101110001110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000001100000000000000000000000000000000000000000000000011100000000000000111111111111111111111111111110111110111110000000111111111111110001111011000011111111111001111111111011101111101110001111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000111000000000000000000000000000000000000000000000000111000000000000111111111111111111111111111110111110111110000000111111111111110001110011001001111111100011111111111011011111101110011111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000111000000000000000000000000000000000000000000000011100000000000111111111111111111111111111111111110111110000001111111111111110001110111001100111111001111111111110111011111101110011111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000001110000000000000000000000000000000000000000000001111000000000111111111111111111111111111101111101111110000001111111111111110001100111011110011100011111111111110110111111101100011111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000011100000000000000000000000000000000000000000000011100000000111111111111111111111111111101111101111110000001111111111111110011101111011111001001111111111111101110111111101100000111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000011000000000000000000000000000000000000000000001110000000111111111111111111111111111101111101111100000001111111111111110011001111011111100011111111111111101101111111101100000011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000110000000000000000000000000000000000000000000011100000111111111111111111111111111111111101111100000001111111111111110011011111011111000111111111111111001101111111101100000011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000001100000000000000000000000000000000000000000001110000111111111111111111111111111011111011111100000001111111111111110010011111011100011011111111111111011011111111101111110011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000001000000000000000000000000000000000000000000011000111111111111111111111111111011111011111000000011011111111111110010111111011001111101111111111110010011111111101001110011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000010000000000000000000000000000010000000000000000000000000000000000000000001010111111111111111111111111111111111011111000000011001111111111110000111100000111111100111111111110110111111111100001110011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110111111111111000000011001111111111110001110000000111111110111111111100101111111110000111110011000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110111110111111000000011001111111111110001100000000001111111011111111101001111111001100111110000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000001100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110111110111110000000011001111111111110011000000000000111111101111111011011111100111110111110001110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000100000001000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110111110000000011001111111111100010000100000000011111111111111010111110011111110111110111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000011001111111111100100001100000000000101111111110101111001111111110111110111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111101111101111110000000110001111111111101000011110000011000010111111110011100111111111110111110111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111101111101111100000000110001111111111101000111110000001100001111111100011011111111111110111100111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111101000000110001111111111101000111110000001110001111111101111111111111111110111101111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000001000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111111111111101000000110001111111111101001111110000111111001111111111111111011111111110111101111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000001000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111011111111111011000000110001111111111101001110000000111111101111111111111110110000111110111101111100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111011111111111011000000100000111111111101001100010000111111101111111111111110000000011110011101111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000001101111111111111111111111111011111111111011100000100000111111111101001100010000001111111111111111111000000000001110011001111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000010000000000000000000000000000000000000000000000000000000000000000000000001101111111111111111111111111111111111111111100000100000111111111101111100000000001111111111111111110000000110001110011011111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000010000000000000000000000000000000000000000000000000000000000000000000000001101111111111111111111111110111111111110111100000100000111111111101111100000000011111111111111111111000000011000111011011111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000001101111111111111111111111110111111111110111100000100000111111111101111100000000011111111111111111111110000011100111010011111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000001000000000000000000000000000000000000000000000000000000000000001101111111111111111111111110111111111110111110000100000111111111011111100000000011111111111111111111111000011100111010111111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000001100000000000000000000000000000000000000000000000000000000011101111111111111111111111111111111111101111110000000010111111111011111100000000011111111111111111111111000111100011010111111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11001111111111100000000000100000000000000000000000000000000000000000000000000000011101111111111111111111111111111111111101111110000000010011111111011111100000000011111111111111111111110001111110011000111111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000111111111111111000000000110000000000000000000000000000000000000000000000000011101111111111111111111111101111111111101111111000000110011111111011111100000000011111111111111111111000011111110011000111111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000110111111111111000000000010000000000000000000000000000000000000000000000011101111111111111111111111101111111111101111111000000110011111111011111101000000111111111111111111111001001111110011001111111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000001111111111111100000000001000000000000000000000000000000000000000000011101111111111111111111111101111111111011111111100000101011111111011111101000110111111111111111111110000000011110010001111111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000111111111111110000000000000000000000000000000000000000000000000111101000111111111111111111111111111111011111111100000101011111111011111101101110111111111111111111110000000111110010001111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000001111111111111000000000000000000000000000000000000000000000111000110001111111111111111011111111111011111111100000111011111111011111101111101111111111111111111110000000111110010001111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000011111111111100000000000000000000000000000000000000000111001111110011111111111111011111111111011111111110000111011111111011111100111111111111111111111111110000000111110100001111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11001000000000000000000000000000111111111110000000000000000000000000000000000000111011111111000000011111111011111111110111111111110000111011111111011111110111011111111111111111111110000000111100100011111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11001111100000000000000000000000000001111111111000000000000000000000000000000001110011111111111111001111111011111111110111111111110000111101111111011111110000111111111111111111111100000000111100100011111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10001011111111110000000000000000000000000111111111100000000000000000000000000001110111111111111111110111111111111111110111111111110000111101111111011111111001111111111111111111111100000001111111000011111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000100011111111100000000000000000000000001111111100000000000000000000000001100111111111111111110011110111111111110111111111110100111101111111111111111111111111111111111111111100000001111111000011111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000011111111110000000000000000000000000011111110000000000000000000001101111111111111111111011110111111111101111111111110110111101111111111111111111111111111111111111111100001001111110000011111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000011111111100000000000000000000000001111111000000000000000001001111111111111111111001110111111111101111111111110110111101111111111111111111111111111111111111111100111011111110000011111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000111100000000000000000000000000001111000000000000000011111111111111111111101110111111111101111111111110110111101111111111111111111111111111111111111111100111011111100000111111100000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000111000000000000011111111111111111111101111111111111101111111111110111011110111111111111111111111111111111111111111110111111111100000111111100000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111100111111111111111111111111110111011110111111111111111111111111111111111111111110000111111100000111111100000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000100111111111011111111111110001111111111011111111111110111011110111111111111111111111111111111111111111111001111111010000111111100000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000100111111111011111111111110100111111111011111111111110011101110111111111111111111111111111111111111111111111111111010001111111000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000101111111110011111111111110110011111111011111111111111011100111011111011111111111111111111111111111111111111111110010001111111000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111110111100111111011111111111111111110011011111011111111111111111111111111111111111111111110110001111111000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111111111110111111001110111111111111111111111000011111011111111111111111111111111111111111111111110100001111110000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000111111111111111111100110111111111111111111111110011111011111111111111111111111111111111111111111110100001111110000010011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000011111111111011111111000111111111111111111111111111111011111111111111111111111111111111111111111110010011111100000010011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000111101111000000000111111111011111111100111111111111111111111111101111011111111111111111111111111111111111111111110010011111101100011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11001100000000000000000000000000000000000000000000000000000000000000000000000111001110000000000001111111011111111110011111111111111111111111101111001111111111111111111111111111111111111111110110011111101100011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000100100011000000000000000000000000000000000000000000000000000000000000000010011000000000000000111111011111111111101111111111111111111111101111001111111111111111111111111111111111111111110110011111011100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000001111011111111111110011111111111111111111101111010111111111111111111111111111111111111111110110111111011000111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000111101111111111111001111111111111111111110111010011111111111111111111111111111111111111110110111110011000111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001101111111111111100111111111111111111110111011011111111111111111110000011111111111111110110111110111000111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110111111111111111111110111011001111111111111111111111001111111111111111110111110111000111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111011111111111111111110111011110111111111111111111111111111111111111101100111101111001011100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000000000000111111111111111011111111111111111111011011111011111111111111111111111111111111111101101111101111011011100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000000000111111111111111101111111111111111111011010111001111111111111111111111111111111111011101111011110011011110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110001000000000000011111111111111100011111111111111111011010111100111111111111111111111111111111111011101111011110011011110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000010001101111111111111111111010010000000000000000000000000000000000000000000111111110011100000000000011111111111111110000110000000000001101010111111011111111111111111111111111111110111101110111110111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100010010011111111111111111111111111111111111111111111111111111111110000000000000111111110011100000000000011111111111111110000111110011111100001010111111101111111111111111111111111111101111101110111110111101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100010110111111111111111111111111111111111111111111111111111111111100000000000001111111110111100000000000011111111111111110000011111001111111001000111111100111111111111111111111111111001111101101111100111101110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100010111001111111111111111111111111111111111111111111111111110000000000000000001111111100111101000000000011111111111111111000001111110111111101101111111111011111111111111111111111110011111011001111101111100111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111100100000000011111111111111111010000111111001111110101111111111100111111111111111111111001111111011011111111111110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111101110000000011111111111111111011000111111100111110001111111111110011111111111111111110011111111010111111111111110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001110000000011111111111111111101100011111110011110001111111111111000111111111111110001111111111010111111111111110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111011110000000011111111111111111111100011111111001111001111111111111110011111111111000111111111111001111111111111110011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111011100000000011111111111111111111110001111111100111001111111111111111100111110000111111111111110011111111111111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111001110100000000000000000000000000000000000000000000000000000000000000000000111111110111111011100000000011111111111111111111110001111111100011101111111111111111100000000111111111111111110011111111111111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000100000000000000000000000000000000000000000000000000000000000000000000000111111110111111011100000000011111111111111111111110001111111111001100111111111111111101111111111111111111111110111111111111111111001101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000101111111101111111111100000000011111111111111111111111000111111110100100011111111111111101111111111111111111111111111111111111111111101101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000001111111111101111110111100000001011111111111111111111111000111111110110010001111111111111101111111111111111111111111111111111111111111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000001111111111101111110111100000001011111111111111111111111100111111110111010000111111111111111111111111111111111111111111111111111111111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000011111111111001111110111100000011011111111111111111111111100111111111111110000011111111111011111111111111111111111111111111111111111111100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000011111111111011111110111100000110111111111111111111111111100011111111011111000001111111111011111111111111111111111111111111111111111111110111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000111111111111011111110111000000110111111111111111111111111100011111111011111000000111111111011111111111111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000000111111111110011111101111011111101111111111111111111111111100011111111011111101000111111111011111111111111111111111111111111111111111111110011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000001111111111110111111101111011111001111111111111111111111111100011111111011111101100011111111011111111111111111111111111111111111111111111111011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000001111111111100111111101111011111011111111111111111111111111100011111111011111100100001111111011111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000011111111111001111111011111011110111111111111111111111111111100001111111111111110110000111111001111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000011111110000011111111011110111100111111111111111111111111111110001111111101111110011000011111101111111111111111111111111111111111111111111111001101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000000000000011111111110111110111001111111111111111111111111111110001111101101111111011100011111100111111111111111111111111111111111111111111111101101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000000110111111111111111001111101110010111111111111111111111111111100001111101111111111011100001111110000001111111111111111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000001110111111111111110011111101110110011111111111111111111111111100001111101111111111001110000001110000000011111111111111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000001111011111111111000111111011101111001111111111111111111111111100001111101111111111101111000000110000000001111111111111111111111111111111111111100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000011111001111111110011111110111001111101111111111111111111111111100001111110111111111100111000010011000000000111111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000000000000000000000000000000000000000000000000011111101111111000111111100110011111110111111111111111111111111000000111110111111111110111100001001010000000011111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000000000000000000000000000000000000000000000000111111110111100101111111001101011111111011111111111111111111111000000111110111111111110111110000101111110000001111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111110000000000000000000000000000000000000000000000000000000111111111000001110111110010011011111111100111111111111111111110000000111110111111111110011110000100111111100000011111111111111111111111111111111111011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111110000000000000000000000000000000000000000000000000000001111111111100111110011100100111011111111100000111111111111111110000110111110111111111111011111000011111111100001000111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111000000000000000000000000000000000000000000000000000001111111111111111111100000011111111111111101100000001111111111100000110111110111111111111011111100001111111110000110001111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111110111111111101110000000001111111000001110111110111111111111001111100000111111110000111110011111111111111111111111111111001101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111110111111111101110000001000111110000011110111110111111111111101111110000011111110000111111001111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111110111111111101110000001111111100000011110111110111111111111101111110000011111110000111111100111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110111111111101110000001111111000000111110111110111111111111101111111000001111110000111111110111111111111111111111111111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111000000000000000000000000000000000000000000000001111111111111111111111111111111101111111111101110000000111110000001111110111110111111111111110111111100000011110000111111111011111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111101111111111111111010000111100000011111110111110111111111111110111111110000000000000011111111011111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111111101111111111111111010000010000000111111110111110111111111111110011111111000000000000011111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111100000000000000000000000000000000000000000111111111111111111111111111111111101111111111011111011000000000001111111110111110111111111111111011111111100000000000011111111101111111111111111111111111110011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111101111111111011111011100000000001111111110111110011111111111111011111111110000000000111111111101111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111111011111111111011111011111000000011111111110111110011111111111111011111111111000000000111111111101111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111100000000000000000000000000000000000111111111111111111111111111111111111011111111111011111001111111000111111111110111110011111111111111101111111110110000000111111111111111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111011111111111011111101111111111111111111110111111011111111111111101111111111011000000111111111110111111111111111111111111111001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111100000000000000000000000000000011111111111111111111111111111111111111011111111111011111101111111111111111111110111111011111111111111111111111111101100001111111111110111111111111111111111111111101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111011111100111111111111111111110111111011111111111111111111111111100111111111111111110111111111111111111111111111101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111110111111111110011111110111111111111111111110111111011111111111111111111111111110111111111111111011111111111111111111111111111101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111110111111111110111111110011111111111111111110111110011111111111111111111111111111011111111111111100111111111111111111111111111110111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111110111111111110111111111011111111111111111110111110011111111111111111111111111111101111111111111110011111111111111111111111111110111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111110111111111110111111111101111111111111111110111110001111111111111111111111111111110111111111111111011111111111111111111111111110111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111110111111111110011111111111111111111100101111111111111111111111111111110111111111111111001111111111111111111111111110011101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111101111111111110111111111111001111111111111111111101101111111111111111111111111111111011111111111111101111111111111111111111111111011101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110111111111111000011111111111111111101101111111111111111111111111111111101111111111111110111111111111111111111111111011111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110111111111111010000000001111111111001101111111111111111111111111111111101111111111111110111111111111111111111111111011111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110111111111111101110000111111111111011101111111111111111111111111111111110111111111111111011111111111111111111111111001110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111111111101111111111111111110011101111111111111111111111111111111110111111111111111011111111111111111111111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111111111100111111111111111110111101111111111111111111111111111111110111111111111111101111111111111111111111111101111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111101111111111111110111111111111111100111100111111111111111111111111111111111011111111111111101111111111111111111111111101111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111101111111111111110111111111111111101111110111111111111111111111111111111111011111111111111110111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111101111111111111111011111111111111001111110111111111111111111111111111111111011111111111111110111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111111111111111011111111111111011111110111111111111111111111111111111111011111111111111111011111111111111111111111110111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111111111111111001111111111110011111110111111111111111111111111111111111011111111111111111011111111111111111111111110111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111111111111111101111111111110111111110111111111111111111111111111111111011111111111111111011111111111111111111111110111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111111111111111101111111111100111111110111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111111111111111100111111111111111111110111111111111111111111111111111111111111111111111111101111111111111111111111111011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111100111111111111111111110111111111111111111111111111111111101111111111111111101111111111111111111111111011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111100011111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111101111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111001111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111101111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111011111111111111111111111111111111111111111011111111111111111111111111111111101111111111111111101111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111011111111111111111110111111111111111111111011111111111111111111111111111111101111111111111111101111111111111111111111111101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111110111111111111111111111011111111111111111111111111111111101111111111111111101111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111111111111111011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111111111111111011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111101001111111111111111111111111111111111111111111111011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111011111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111001111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111110111111111111111111111101111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111110111111111111111111111101111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111101111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111101111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111100111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111011111111111111111111111111111110111111011111011111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111011111111111111111111111111111110111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111110111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111110111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111110011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111110111111111111111111111111011111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111011111101111101111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111110111111111111111111111111011111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111011111101111110111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111110111111111111111111111111011111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111110111111111111111111111111011111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111110111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111110111111111111111111111111111111111101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111110111111111111111111111111101111111111111111111111111111111111111111111001111111111111111111110111111111111111111111111111111111101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111110111111111111111111111111111111111101111110111111011111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111110111111111111111111111111111111111101111111111111011111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111110111111111111111111111111111111111101111111011111011111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110111111111111111111111111110111111111111111111111111111111111111111110011111111111111111111110111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110111111111111111111111111110111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111011111101111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100111111110111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100111111110111111111111111111111111111011111111111111111111111111111111111111101111111111111111111111101111111111111111111111111111111111110111111101111101111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100111111110111111111111111111111111111011111111111111111111111111111111111111001111111111110111111111101111111111111111111111111111111111110111111101111110111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111011111111111111111111111111111111111111001111111111110111111111101111111111111111111111111111111111111011111111111110111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111110111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111110111110111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111001111110111111011111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111101111111111111011111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101111111011111011111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111011111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111101111111111111011111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111011111111111111111111111111111111111111111111111110011111110111111111111111111111111111111111111111101111111111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110111111111111111111111111111111111111111100111111111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111101111111111111111111111111111111111111111111111110011111110011111111111111111111111111111111111111100111111111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111110111111111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111110111111111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111101111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111");
BEGIN 
	--WRITE PROCESS
		
   read_process: PROCESS(clk)
	BEGIN 
	   IF (rising_edge(clk)) THEN
				data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;