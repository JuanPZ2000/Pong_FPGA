LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY romGreen IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=320;
					ADDR_WIDTH	:	INTEGER:=8);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF romGreen IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111100000000011111111111111111111000000111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100","11111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000011111111111111111000111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000","11111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000011111111111111100011111111111111111111110000000011100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000","11111111111111111111111111100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000001111111111110011111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000","11111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000111111111001111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000","11111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000","11111111111111111111111110011100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000","11111111111111111111111100001100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111100000000011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000","11111111111111111111111000001111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000011100111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000","11111111111111111111111000000011100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111000000000011011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000","11111111111111111111110000000001100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111100000000010111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000","11111111111111111111100000000000001100000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111110111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000","11111111111111111111000000000000001110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000001111101111111111111111111111111111111111111111111111111110111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111111110000010000000000111000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000011111001111111111111111111111111111111111111111111111111110111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111111110000000000000000011110000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000111111011111111111111111111111111111111111111111111111111111011111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111111100000000000000000000111000000000000000000000000000000000000000111111111111111111111111111111111111111111111101110000000101110011111111111111111111111111111111111111111111111111111001111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000","11111111111111111000000000000000000000011100000000000000000000000000000000000000111111111111111111111111111111111111111111111011111110000000000011111111111111111111111111111111111111111111111111111001111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111011111111000000000101111111111111111111111101111111111111111111111111111000111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111111000000000000001000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111110111001111000000000100000000000011101111111001111111111111111111111111111001011100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111110000000000000000110000000000000000000000000000000000000000000000011111111111111111111111111111111111111111110111000111000000000000000000000000000001111011111111111111111111111111111101001110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000","11111111111111110000000000000000001000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000010000000000000000000000000000000010000011111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000","11111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111101110000000000000000000000000000000000000000000000011111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000","11111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111101110000000000000000000000000000000000000000000000000000011111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111111000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111011100000000000000000000000000000000000000000000000000000000000111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000","11111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111011100000000000000000000000000000000000000000000000000000000000001111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000101111","11111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000110001111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111","11111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111110111100000000000000000000000000000000000000000000000000000000000000000001111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111","11111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111110111000000000000000000000000000000000000000000000000000000000000000000001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000001000100000000000000000000000000000000000000000000000000000000100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111101111000110000000000011000100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111101111000110000000000011000100000000000100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111011110001110000000000111001100000000010100000000010000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111011110001110000000000111001000000000111111000000110000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111011110001110000000001111011100000000111110000000111000011000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110111110011110000000001111111110000000111110000001111111111111000000000100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110111100011110000000011111111110000001111110000001111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110111100011100000000111111111110000001111110000011111111111111110000010000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111100111100000000111111111110000011111100000111111111111111100000100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111101111100111100000001111111111110000011111100000111111111111111000000000001000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111101111000111100000001111111111110000011111000000111111111111011000000000011001000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111101111001111000000001111111111110000111100000001111111111111110001000000011001000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111011111001111000000011111111111110000111100000001111111111111100000000000110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111011111001111000000011111111111110000111100000001111111111101000000000100110010000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111011110001111000000011111111111110000111100000011111111111110000000000001110100001100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110011110000000111111111111110001111001000011111111111100000000001001100100001110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110111110011110000000111111111111100001110001000001111111110001000000000001001100001110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110111100011110000000111111111111100001110011000001111111100010000000010011001110001100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110111100011110000000111111111111100001100111000100111110000100000001110010011110001100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111101111100111100000000111111111111100001100111001110011100000000000111110110011110001100001000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111101111100111100000001111111111111100001001111001111000000100001111111100100111110001100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111101111100111100000001111111111111100001001111011111100000001111111111101100111110001000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011111001111100000001111111111111100001011111011110000011111111111111001001111110000100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011111001111000000001001111111111100010011110011100011011111111111111011011111111001111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011111001111000000001001111111111100010111110010001111001111111111110010011111111000001100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110011111000000001001111111111100000111100000011111100111111111110100111111111000001110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110111110011111000000011001111111111100001110000000111111110111111111100100111111110000110110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110111110011110000000011001111111111100001100000000001111111011111111101001111111000100101110000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110111110011110000000011001111111111100011000000000000111111101111111000011111100011100111110000100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110111100111110000000011001111111111100000000000000000001101101111111000111110001111100111110011100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101111100111100000000010001111111111100100001100000000000100111111110000111000111111100111100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101111100111100000000010001111111111100000011110000001000000111111100001100011111111100111100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101111101111100000000010001111111111100000111110000001100000111111100011001111111111100111100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101111001111101000000010000111111111101000111110000001110001111111001111111111111111100011100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111001111001000000100000111111111101001111100000001111001111111111111110011111111100011100111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011111001111011000000100000111111111101001100000000111111101111111111111100100000111110011001111100010011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011111011111011000000100000111111111101001100000000111111101111111111111110000000011110011001111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011111011111011100000100000111111111001001100000000001111111111111111111000000000001110011001111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110011110011100000100000111111111001001100000000001111111111111111110000000110001110011001111100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111110011110111100000100000111111111001111100000000001111111111111111110000000011000110010011111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111110111110111100000000000111111111001111100000000011111111111111111111110000011000110010011111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111110111100111110000000000011111111001111100000000011111111111111111111111000011100010010011111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111110111101111110000000010011111111011111100000000011111111111111111111111000011100011000111111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111101111101111110000000010011111111011111100000000011111111111111111111110001111110011000111111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000110011110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111101111101111111000000010010111111011111100000000011111111111111111111000001111110011000111111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000001111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111101111001111111000000100011111111011111100000000111111111111111111110000000111110000000111111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000011000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111101111001111111100000100011111111011111100000100111111111111111111110000000011110000000111111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111101111011111111100000100011111111011111100000100111111111111111111110000000011110010000111111000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001111111111111111011111011111011111111100000100010111111011111100001101111111111111111111110000000111110000000111111000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100011111111111111011111011110011111111100000110001111111011111100001101111111111111111111110000000111110000000111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11001000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000011111111011111011110011111111110000110001111110011111110000011111111111111111111100000000111100100001111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11001111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111011111111110111111111110000110001111110011111110000011111111111111111111100000000111100000001111111000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000011100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100111111111111111110111111111110000110001111110011111110000111111111111111111111100000001111111000001111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110011110111111111100111111111110100110001111110011111111111111111111111111111111100000001111111000001111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011110111111110101111111111110110111000111110011111111111111111111111111111111100001001111110000001111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111001110111111111101111111111110110111000111110011111111111111111111111111111111100001011111110000011111110000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111101110111111111101111111111110110111100111110011111111111111111111111111111111100001011111100000011111100000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100001111111101110111111111001111111111110111011100111110011111111011111111111111111111111110010111111100000011111100000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000011111100111111111111001111111111110111011110111110011111100001111111111111111111111110000111111000000011111100000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000011111100001111111111011111111111110011011110011110011111000001111111111111111111110110001111111000000111111000000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111110100111111111011111111111110011101110011110011111000001111111111111111111111111111111111010000111111000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111110110001111110011111111111111011100110011110011111100001111111111111111111111111111111110000000111111000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000001111101110010000001111110111100111110011111111111111111110011011110011111110011111111111111111111111111111111110000000111110000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000011111001100001000001111110111110001110111111111111111111111000011110001111111111111111111111111111111111111111110100000111110000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000010000111110011111100010111111111111111111111110001110001111111111111111111111111111111111111111100000001111010000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000011100001000000001000111111011111110000111111111111111111111111001110010111111111111111111111111111111111100011110010001111100000010001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000011100010000000000010111111011111111100111111111111111111111111101110000111111111111111111111111111111111100001110010001111101100010001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000011000100000000000000111111011111111110011111111111111111111111101110001011111111111111111111111111111111110001110110011111001100010001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000011111011111111111101111111111111111111111100110000011111111111111111111111111111111101001100110011111001100010001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111001111111111110011111111111111111111100110010001111111111111111111111111111111111111100110011111011000110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001111111111111001111111111111111111110110010001111111111111111111111111111111111111100110011110011000111001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111111111111100111111111111111111110110011001111111111111111110000011111111111111100110111110111000111000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110111111111111111111110010011000111111111111111111111001111111111111100110111100111000011000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111011111111111111111110011011000011111111111111111111111111111111111101100111101111001011000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111111111111111011111111111111111111011010010011111111111111111111111111111111111001100111001111011011100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","10000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000000000111111111111111101111111111111111111011010001001111111111111111111111111111111111011100111011110011001100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110001000000000000011111111111111100011111111111111111001010000100111111111111111111111111111111110011101110011110011001100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110011100000000000011111111111111110000110000000000001101010000010011111111111111111111111111111110111101110111110111101100011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000010000000000000000000000000000000000000000000000000000000000000000000000000111111110011100000000000011111111111111110000111110011111100001010000001001111111111111111111111111111101111101100111110111101110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100010000000000000000000000000000000000000000000000000000000000000000000000000000111111100011100000000000011111111111111110000011111001111111001000000000100111111111111111111111111111001111101101111100111100110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100010000000000000000000000000000000000000000000000000000000000000000000000000001111111100111100000000000011111111111111111000001111110111111100000000000010001111111111111111111111110011111001001111101111100110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111100000000000011111111111111111010000111111001111110000000000001000111111111111111111111001111111001011111111111110110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111000110000000011111111111111111001000111111100111110000000000000100011111111111111111100011111111010011111111111110010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11100000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111001110000000011111111111111111101100011111110011110000000000000000000111111111111110001111111111000111111111111110010001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111001100000000011111111111111111111100011111111001111000000000000000100001111111110000111111111110001111111111111110011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11110000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111011100000000011111111111111111111110001111111100111000000000000000000000111100000111111111111110011111111111111111011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111011100000000001111111111111111111110001111111100011100100000000000000100000000111111111111111110011111111111111111001001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111011100000000001111111111111111111110001111111111001100000000000000000001111111111111111111111110111111111111111111001000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000100111111100111110011100000000001111111111111111111111000111111110100100000000000000000001111111111111111111111111111111111111111111101100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000000000111111101111110111100000000000001111111111111111111000111111110110010000000000000000001111111111111111111111111111111111111111111101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111000000000000000000000000000000000000000000000000000000000000000000000001000111111101111110111100000000000000011111111111111111000111111110111010000000000000000011111111111111111111111111111111111111111111100100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000011111001111110111100000000010000011111111111111111100111111111111110000000000000000011111111111111111111111111111111111111111111100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000010000001111001111110111000000010000000001111111111111111100011111111111111000000000000000011111111111111111111111111111111111111111111110110011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111100000000000000000000000000000000000000000000000000000000000000000000000000000111011111100111000000100100000000111111111111111100011111111011111000000100000000011111111111111111111111111111111111111111111110110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000000000000000010011111100111001001000000000000111111111111111100011111111011111101000000000000011111111111111111111111111111111111111111111110010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111110000000000000000000000000000000000000000000000000000000000000000000000000000010010000000111000000001000000000011111111111111100011111111011111101100000000000011111111111111111111111111111111111111111111111011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000001000000000100100000000011000000010000000000001111111111111100011111111011111100100000000000011111111111111111111111111111111111111111111111011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111000000000000000000000000000000000000000000000000000000000000000000011001100000000001001010000000000000000000000111111111111100001111111111111110110000100000001111111111111111111111111111111111111111111111001001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000111111111111000001111111101111110011000010000001111111111111111111111111111111111111111111111001001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000000000000000000010100000000001000100000000000000011111111111000001111111101111111011100001000000111111111111111111111111111111111111111111111101101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111100000000000000000000000000000000000000000000000000000000000000110000000000000011000000000100010000000000000000001111111110000001111101111111111011100000110000000001111111111111111111111111111111111111111101100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111110000000000000000000000000000000000000000000000000000000000001110000000000000100001001001100110000000000000000001111111110100001111101111111111001110000000100000000011111111111111111111111111111111111111100100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000001111000000000000000010010001001111001000000000000000111111100100001111101111111111101111000000010000000001111111111111111111111111111111111111100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000011111000000000100000000000010001110100100000000000000111111000000001111110111111111100111000000010000000000111111111111111111111111111111111111110110111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111000000000000000000000000000000000000000000000000000000000011111100000010000100000000100011110100000000000000000011110001000000111110111111111110111100000001000000000011111111111111111111111111111111111110110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111100000000000000000000000000000000000000000000000000000000111111110011000000100000001001011110110001000000000000001100000000000111110111111111110111110000000100000000001111111111111111111111111111111111110010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111110000000000000000000000000000000000000000000000000000000111111111000001110000000010011011100111000001100000000000000010000000111110111111111110011110000000100011100000011111111111111111111111111111111111011011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111110000000000000000000000000000000000000000000000000000001111111111100111110001100000111011100111100000000110000000000100000110111110111111111111011111000000000011100001000111111111111111111111111111111111011011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111000000000000000000000000000000000000000000000000000001111111111111111111100000011111011101111101100000000000000000100000110111110111111111111011111100000000111110000110001111111111111111111111111111111001001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111110111101111101110000000000000001000001110111110111111111111001111100000101111110000111110011111111111111111111111111111001001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111110111101111101110000000000000010000011110111110111111111111101111110000011111110000111111001111111111111111111111111111101101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111110111001111101110000001111000100000011110111110111111111111101111110000001111110000111111100111111111111111111111111111101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111110111001111001110000000000001000000111110111110111111111111101111111000000111110000111111110111111111111111111111111111100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111000000000000000000000000000000000000000000000001111111111111111111111111111111101111011111001110000000100110000001111110111110111111111111110111111100000011110000111111111011111111111111111111111111100110111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111101111011111001111010000001000000011111110111110111111111111110111111110000000000000011111111011111111111111111111111111110110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111111101111011111011111010000000000000111111110111110111111111111111011111111000000000000011111111111111111111111111111111111110010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111101110011111011111011000000000000111111110111110011111111111111011111111100000000000011111111101111111111111111111111111110011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111100000000000000000000000000000000000000001111111111111111111111111111111111101110011111011111011100000000001111111110111110011111111111111011111111110000000000111111111101111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111110000000000000000000000000000000000000011111111111111111111111111111111111011110111111011111011111000000011111111110111110011111111111111011111111111000000000111111111101111111111111111111111111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111100000000000000000000000000000000000111111111111111111111111111111111111011110111111011111001111111000111111111110111110011111111111111101111111110110000000111111111111111111111111111111111111111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111011110111111011111101111111111111111111110111111011111111111111101111111111011000000111111111110111111111111111111111111111001100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111000000000000000000000000000000011111111111111111111111111111111111111011110111110011111101111111111111111111110111111011111111111111111111111111101100001111111111110111111111111111111111111111101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111011100111110011111100111111111111111111110111111011111111111111111111111111100111111111111111110111111111111111111111111111101100111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111110111100111110011111110111111111111111111110111111011111111111111111111111111110111111111111111011111111111111111111111111111100110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111110111100111110111111110011111111111111111110111110011111111111111111111111111111011111111111111100111111111111111111111111111100110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111110111101111110111111111001111111111111111110111110011111111111111111111111111111101111111111111110011111111111111111111111111110110011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111110111101111110111111111101111111111111111110111110001111111111111111111111111111110111111111111111011111111111111111111111111110011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111101111101111110111111111110011111111111111111111100101111111111111111111111111111110111111111111111001111111111111111111111111110011001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111101111101111110111111111111001111111111111111111101101111111111111111111111111111111011111111111111101111111111111111111111111111011001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111110111111111111000011111111111111111101101111111111111111111111111111111101111111111111110111111111111111111111111111011100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111001111100111111111111010000000001111111111011101111111111111111111111111111111101111111111111110111111111111111111111111111001100111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111001111100111111100000000000000000111111110000000000111111111111111110000000000000011110000000000011111000000000011111111111001110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111100111111100000000000000000001111110000000000111111111111111100000000000000011110000000000011111000000000011111111111101110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111100111111100000000000000000000111110000000000111111111111111100000000000000001110000000000001110000000000011111111111101110011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111101111111100000000000000000000011100000000000111111111111111100000000000000001111000000000001110000000000111111111111100110011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111101111111100000000000000000000001100000000000111111111111111100000000000000001111000000000000100000000000111111111111100111011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111","01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111101111111100000000000000000000001000000000000111111111111111000000000000000001111100000000000100000000001111111111111110111001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111","01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110011111101111111100000000000000000000000010000000000111111111111111000000000000000000111110000000000000000000001111111111111110111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110011111101111111100000000000100000000000010000000000111111111111111000000000000000000111110000000000000000000011111111111111110111101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110011111101111111100000000001110000000000110000000000111111111111111000000000000000000111110000000000000000000011111111111111110011100111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110011111101111111100000000000110000000000110000000000111111111111110000000000000000000111111000000000000000000111111111111111111011110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111111101111111100000000000110000000000110000000000111111111111110000000000000000000011111100000000000000000111111111111111111011111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110111111001111111100000000000110000000000110000000000111111111111110000000000000000000011111100000000000000001111111111111111111011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111101111111100000000000010000000000110000000000111111111111110000000000000000000011111110000000000000001111111111111111111001111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111111111111100000000000000000000000110000000000111111111111100000000001000000000011111110000000000000011111111111111111111001111011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111011111111100000000000000000000000110000000000111111111111100000000001100000000001111111000000000000011111111111111111111101111001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111100111111011111111100000000000000000000001110000000000111111111111100000000001100000000001111111000000000000111111111111111111111101111001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111111011111111100000000000000000000001110000000000111111111111000000000001100000000001111111100000000000111111111111111111111100111101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111100000000000000000000011110000000000111111111111000000000011100000000001111111100000000001111111111111111111111100111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111100000000000000000000011110000000000111111111111000000000000000000000000111111100000000001111111111111111111111110111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101111111011111111100000000000000000000111110000000000111111111111000000000000000000000000111111100000000001111111111111111111111110111110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101111011011111111100000000000100000011111110000000000111111111110000000000000000000000000111111100000000001111111111111111111111110111110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110011111111100000000000111111111111110000000000111111111110000000000000000000000000011111100000000001111111111111111111111110011110011110111111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110011111111100000000000011111111111110000000000111111111110000000000000000000000000011111100000000001111111111111111111111110011110011111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110011111111100000000000011111111111110000000000000000000110000000000000000000000000011111100000000001111111111111111111111111011111011111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100000000001011111111111110000000000000000000100000000000000000000000000011111100000000001111111111111111111111111011111001111011111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111111100000000001011111111111110000000000000000000100000000000000000000000000001111100000000001111111111111111111111111011111001111101111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111111100000000001011111111111110000000000000000000100000000001111111100000000001111100000000001111111111111111111111111001111001111101111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111111100000000001011111111111110000000000000000000100000000001111111100000000001111100000000001111111111111111111111111001111101111101111111111111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111110111111111100000000001101111111111110000000000000000000000000000001111111100000000000111100000000001111111111111111111111111101111100111110111111111111111111111111111111111111111111111111111111111111111111111111111111","01111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111001111110111111111100000000001101111111111110000000000000000000000000000011111111100000000000111100000000001111111111111111111111111101111110111110111111111111111111111111111111111111111111111111111111111111111111111111111111","01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111111110000000001101111111111111000000000000000000000000000011111111000000000000111100000000001111111111111111111111111101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111","11101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111100111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111","00000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111110111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111100111110111111011111111111111111111111111111111111111111111111111111111111111111111111111111","00000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111011111111111111111111111111111110111110011111011111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111011111111111111111111111111111110111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111","00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111110011111011111101111111111111111111111111111111111111111111111111111111111111111111111111111","11111001110101111111111111111111111111111111111111111111111111111111111111111111111111101111110011111100111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111110011111001111101111111111111111111111111111111111111111111111111111111111111111111111111111","00000100000111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111100111111111111111111111111011111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111011111001111101111111111111111111111111111111111111111111111111111111111111111111111111111","00000000101111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111110111111111111111111111111011111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111011111101111110111111111111111111111111111111111111111111111111111111111111111111111111111","00000000111111111111111111111111111111111111111111111111111111111111111111111111111111101111110011111110111111111111111111111111011111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000001111111111111111111111111111111111111111111111111111111111111111111111111000001101111110011111100111111111111111111111111011111110001111111111111101111011111111111111101111111111111111111111111111111111111111111011111111111001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111","00000111111111111111111111111111111111111111111111111111111111111111111111111111000000101111100011111110111111111111111111111111111111110001111111111111001110011111111111111101111001111111111111111111111111111111100110011111111111101111100111111111111111111111111111111111111111111111111111111111111111111111111111111111","00001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000100001100000100001111100011000000100000011110000011000100110000100001100011000000001110000110001111110000110001100000011000011010000001000100010000111111111111111111111111111111111111111111111111111111111111111111111111111111111","00011111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111000001000000000000011110000001000000100000000001000001000000011100000000000111100000100000100000010000000010000001000100000000011111011111111111111111111111111111111111111111111111111111111111111111111111111","01111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111000000000000000000011110000001000000000000000010000001000000011100001000000111000000000000100000000000100010000000000100000000011111011111111111111111111111111111111111111111111111111111111111111111111111111","11111110111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111100000000100010000011110000000000000110001000010000000000000011100001000000111000010000100100010001000100010001000000100000000011111011111111111111111111111111111111111111111111111111111111111111111111111111","11111100111111111111111111111111111111111111111111111111111111111111111111111110000000100011000000000000100001111000000000100010000111110000000000000100001000010000000000000011100001000000111000010000100100010000000100010001000000100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111","11100110000111111111111111111111111111111111111111111111111111111111111111111110000111000011000000000000110001111001000000100010000111110000001000000110000100000000001000000011100000000000111000000000000100010001000000010001000000000000000011111101111111111111111111111111111111111111111111111111111111111111111111111111","10000000000111111111111111111111111111111111111111111111111111111111111111111110000111000011100000000000000001111000000000100010000111110000001000000110000100001000001000000011110000000000111100000100000100010001000000010001000000000010000001111101111111111111111111111111111111111111111111111111111111111111111111111111","10000000001111111111111111111111111111111111111111111111111111111111111111111111000111000011100000100000100011111100000000100010000111110000011100100111000110001100011000000011110001110001111110000110001100010011100100010001001100100010000001111101111111111111111111111111111111111111111111111111111111111111111111111111","00000000011111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111110111111111111111111111110001011111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111110111111001111101111111111111111111111111111111111111111111111111111111111111111111111111","00000000111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111110111111111111111111111110001011111111111111111111111111111111111111001111111111110111111111101111111111111111111111111111111111110111111001111110111111111111111111111111111111111111111111111111111111111111111111111111","00000001111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111110111111111111111111111111111011111111111111111111111111111111111111001111111111110111111111101111111111111111111111111111111111111011111100111110111111111111111111111111111111111111111111111111111111111111111111111111","00000011110111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111100111110111111111111111111111111111111111111111111111111111111111111111111111111","00000111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111100111110111111111111111111111111111111111111111111111111111111111111111111111111","00001110111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111001111100111110111111111111111111111111111111111111111111111111111111111111111111111111","00110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111001111110111111011111111111111111111111111111111111111111111111111111111111111111111111","00110011111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111001111110011111011111111111111111111111111111111111111111111111111111111111111111111111","10000111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111111111111101111110011111011111111111111111111111111111111111111111111111111111111111111111111111","00111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000011111100111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101111111011111011111111111111111111111111111111111111111111111111111111111111111111111","00111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111011111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111100111111111111011111111111111111111111111111111111111111111111111111111111111111111111","01111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111100111111111111111111111111111111011111111111111111111111111111111111111111111111110011111110111111111111111111111111111111111111111100111011111111001111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111100111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110111111111111111111111111111111111111111100111111111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111100111111111111111111111111111111101111111111111111111111111111111111111111111111110011111110011111111111111111111111111111111111111100111101111111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111110111111011111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111110111101001111101111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111110011101001111100111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111000111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110011111100111110111111111111111111111111111111111111111111111111111111111111111111111");
BEGIN 

	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
		   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;