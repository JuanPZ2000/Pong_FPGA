LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY romBlue2 IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=320;
					ADDR_WIDTH	:	INTEGER:=8);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF romBlue2 IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("00000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000111111110000000000000000000","00000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000001111111100000000000000000000","00000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000011111111000000000000000000000","00000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001110011000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000111111110000000000000000000000","00000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000001110010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001111111100000000000000000000000","00000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000011100000000000000000101111110110000000000000000000000000000000000000000000000000000100000000000000000000000000000000000011111110000000000000000000000000","00000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000011110000000000000000011111100110000000000000000000000000000000000000000000000000001100000000000000000000000000000000000111111100000000000000000000000000","00000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000011100000000000000000111111100100000000000000000000000000000000000000000000000000011000000000000000000000000000000000011111111000000000000000000000000000","00000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011111000000000000001111111101100000000000000000000000000000000000000000000000000110000000000000000000000000000000000111111110000000000000000000000000000","00000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011000000000000000000000000000000001111111001100000000000000000000000000000000000000000000000001110000000000000000000000000000000001111111100000000000000000000000000000","00000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000011100000001111111000000000000000000001111111001100000000000000000000000000000000000000000000000011100000000000000000000000000000000011111111000000000000000000000000000000","00000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000110000111111111111111111110000000000000000111011000000000000000000000000000000000000000000000000011000000000000000000000000000000000111111100000000000000000000000000000000","00000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000001000111111111111111111111110000000011111000111011000000000000000000000000000000000000000000000000110000000000000000000000000000000001111111000000000000000000000000000000000","00000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000011111111111111111111111000011111111111111110110000000000000000000000000000000000000000000000001100000000000000000000000000000000111111110000000000000000000000000000000000","00000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000001111111111111111111111111111111111111111111110110000000000000000000000000010000000000000000000011100000000000000000000000000000001111111100000000000000000000000000000000000","00000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000111000000000000000000011111111111111111111111111111111111111111111111110000000000000000000000000010000000000000000000111000000000000000000000000000000011111111000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000001111100000000000000001111111111111111111111111111111111111111111111111100000000000000000000000011100000000000000000001110000000000000000000000000000000111111100000000000000000000000000000000000000","00000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000111100000000000000011111111111111111111111111111111111111111111111111100000000000000000000000111100000000000000000001110000000000000000000000000000001111111000000100000000000000000000000000000000","00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000111000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000111000000000000000000111100000000000000000000000000000011111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000011000000000000011111111111111111111111111111111111111111111111111111100000000110000000000001110000000000000000001111011000000000000000000000000000111111100000100000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000011000000000000111111111111111111111111111111111111111111111111111111110000001100000000000011110000000000000000011111100000000000000000000000000011111111000001000000000000000000000000000000000000","00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011100000000001111111111111111111111111111111111111111111111111111111110000001110000000000111100000000000000000111111110000000000000000000000000111111110000010000000000000000000000000000000000000","00000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000001111111100000000001110000000001111111111111111111111111111111111111111111111111111111110001111000000000000111100000000000000001111111110000000000000000000000001111111100001100000000000000000000000000000000000000","00000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000001111111110000000011110000000011111011111111111111111111111111111111111111111111111111110000111000000000011111000000000000000011111111100000000000000000000000011111110000011000000000000000000000000000000000000000","00000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000111111011111111111111111111111111111111111111111111111111111011110000000000001111000000000000000111111111000000000000000000000000111111100000100000000000000000000000000000000000000000","00000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000111111111000000001111000001111111011111111111111111111111111111111111111111111111111111001111000000000001111000000000000011111111110000000000000000000000001111111000011000000000000000000000000000000000000000000","00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111110001111110111111111111111111111111111111111111111111111111111111000111000000000001110000000000000111111111110000000000000000000000011111110000110000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000011111111011111100111111111111111111111111101111111111111111111111111111010111000000000001110000000000001111111111100000000000000000000000111111100001100000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000111111111011111100111111111111111111111111101111111111111111111111111111111011100000000001110000000000011111111111000000000000000000000011111111000011000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000111111111011111101111111111111111111111111011111111111111111111111111111111000100000000001110000000000111111111111000000010000000000000111111110001100000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100111111110011111001111111111111111111111110111111111111111111111111111111111100000000000001100000000011111111111110000001100000100000011111111000011100000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111101111111110011111001111111111111111111111110111111111111111111111111111111111100000000000001100000000111111111111110000011100011111110011111110000110000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111110011111011111111111111111111111100111111111111111111111111111111111110000000000001100000011111111111111110000111111111101100111111100011100000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110011110011111111111111111111111101111111111111111111111111111111111110000001111111100000111111111111111100011111111111110111111111000111000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110011110111111111111111011111111001111111111111111111111111111111111111000001111111100111111111111111111011111111111111110111111110001110000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111111100011110111111111111110011111111011111111111111111111111111111111111111000001111111001111111111111111111111111111111111111111111100111100000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111111111100011100111111111111110011111111011111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111110001110000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111111111100011101111111111111110111111110111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111110011100000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110111111111100011101111111111111100111111110111111111111111111111111111101111111111100001111111111111111111111111111111111111111111111111101111000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101111111111100011001111111111111100111111100111111111111111111111111111001111111111110001111111111111111111111111111111111111111111111110011110000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000111101111111111000111001111111111111101111111101111111111111111111111111110011101111111110001111111111111111111111111111111111111111111111100111100000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011101111111111010111011111111111111101111111101111111111111111111111111100011101111111110001111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001011111111111010110011111111111111001111111001111111111111111111111111000011101111111111001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000001011111111111010110011111111111111011111111011111111111111111111111110000111001111111111001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000011111111111010110111111111111111011111111011111111111111111111111100100111001111111111001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000010111111111110010110111111111111111011111110011111111111111111111111000100111001111111111001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100010111111111110110100111111111111110011111110111111111111111111111110000001110001111111111100111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000111111111110110101111111111111110011111110111111111111111111111100000001110001111111111100111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011111111111110001111111111110110001111111111111110111111110111111111111111111111000000011100011111111111100011111111111111111111111111111111111111110000000000000000000000111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000011111111111111101111111111100110001111111111111110111111100111111111111111111110010000011100011111111111101011111111111111111111111111111111111111100000000000000000000011111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000011111111111111001111111111101110011111111111111100111111000111111111111111111100000000011100001111111111100011111111111111111111111111111111111111000000000000000000011111111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000011111111111111001111111111100110011111111111111100111111001111111111111111111001000000111000001111000111110011111111111111111111111111111111111110000000000000000011111111111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000001111111111111011111111111100110011111111111111101111110001111111111111111110010000000111000001111000011110011111111111111111111111111111111111100000000000000111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000001111111111111011111111111000110111111111111111101111110001111111111111111100000000001110000001111000001110001111111111111111111111111111111110000000000000011111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000001111111111111011111111111010110111111111111111101111100000111111111111110000000000001110000011110000000110001111111111111111111111111111111100000000000011111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000001111111111110111111111111010110111111111111111101111001000111111111111100000000000001100100001110000000000001111111111111111111111111111111100000000011111111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000001111111111110111111111111010100111111111111111101111001000011111111111000000000000011101100001110000000000001111111111111111111111111111111000000111111111111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111101111111111110111111111110010100111111111111111101110011001101111111100010000000010011001110001110000000000001111111111111111111111111111111101111111111111111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111101111111111110110101111111111111111001110011011100111111000100000001110111011110001110000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111101111111111110110001111111111111111011100111011110011100000000000111100110011110001100000000001001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111101111111111110110001111111111111111011101111011111001000100000111111101110111110001100000000001001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111111111111111111101111111111100110001111111111111111011001111011111100000000111111111101100111110001100000000001001111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000111111111111111111011111111111101111001111111111111111011011110011111000000111111111111011101111110001100000000001001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011111111111111111011111111111101111011111111111111111011011110011100010011111111111111011011111111001111110000000000111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000111","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000001111111111111111011111111111101111011011111111111111010111110011001111001111111111110011011111111001101110000000000111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111100","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000001111111111111111111111111111001111011011111111111111010111100000011111100111111111110110111111111000011110000000010111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000111110000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000111111111111110111111111111001111011001111111111110001110000000111111110011111111101100111111110000111110000000010111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000111111000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000011111111111110111111111111001111011001111111111110001100000000001111111011111111101101111110000000111110000001010111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011111000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000001111111111110111111111111000110011001111111111110001000000000000111111001111111011011111000011100111110001111010111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011111000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100001111111111110111111111110100110011001111111111110000000000000000001101100111111010111110001111100111110111111010111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111101111111111110100110111001111111111110000001100000000000100111111110100110000111111100111110111111010111111111111111111111111111111111111111111111000000000000000000000000000000000000000011111100000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111101111111111110110110111001111111111110000011110000011000000111111100001100011111111100111110111111010111111111111111111111111111111111111111111110000000000000000000000000000000000000011111100000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111101111111111100010110110001111111111110000111110000001100000111111100011001111111111100111110111111010111111111111111111111111111111111111111111100000000000000000000000000000000000011111110000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100010110110101111111111111000111110000001110001011111000111111111111111100111101111111010111111111111111111111111111111111111111110000000000000000000000000000000000011111110000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111011111111111101010110110101111111111101001111110000111111001111111111111100011111111100111101111111010011111111111111111111111111111111111111100000000000000000000000000000000011111110000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011111111111101010110110101111111111101001110000001111111101111111111111100100000011100111101111111011011111111111111111111111111111111111111100000000000000000000000000000011111111000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011111111111011000010110101111111111101001100010000111111100111111111111110000000011110111101111111011011111111111111111111111111111111111111111000000000000000000000000111111111110000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011111111111011100010100101111111111101001100010000001111111111111111111000000000001110111011111111011011111111111111111111111111111111111111111110000000000000000000111111111111000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111111111111011101010100110111111111101001100000000001111111111111111110000000110001110011011111111011011111111111111111111111111111111111111111111111110000000011111111111111110000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111111111110111101010101100111111111101111100000000011111111111111111110000000011000110011011111111011011111111111111111111111111111111111111111111111111111110111111111111111100000000000000000000000000000000000","11000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111111111110111100000101100111111111101111100000000011111111111111111111110000011000110010011111111011011111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000","11110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111111111110111110100101000111111111101111100000000011111111111111111111111000011100010010111111111011011111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000","00011111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111111111111111110100101010111111111001111100000000011111111111111111111111000111100010010111111111011011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000","00000111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111111111101111110001001010111111111011111100000000011111111111111111111110001111110011000111111111011011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000","00000000010001100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111111111101111111001000010111111111011111100000000011111111111111111111000011111110001001111111111011011111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111111111101111111001000100011111111011111101011010111111111111111111110001001111110000001111111111011011111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101111111111101111111101000100011111111011111101100110111111111111111111110000000011110000001111111111011011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111011111111111011111111100010100011111111011111101111110111111111111111111110000000111110010111111111110011101111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001111111111111111011111111111011111111100000100011111111011111101111111111111111111111111110000000111110010111111111110111101111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111111111111011111111111011111111100000110011111111011111101111111111111111111111111110000000111110001111111111100111101111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000011111111011111111111011111111110000110011111111011111100111011111111111111111111100000000111100101111111111000111101111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000","00001000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111011111111110111111111110000110001111111011111110110111111111111111111111100000000111100001111111111010111101111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100111110111111111110111111111110000110001111111011111111000111111111111111111111100000001111101011111111111010111101111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110011110111111111110111111111110100110001111111011111111111111111111111111111111100000001111111011111111111010111101111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011110111111111111111111111110110111001111111011111111111111111111111111111111100001001111110011111111110010111101111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111001110111111111101111111111110110111001111111011111111111111111111111111111111101111011111110011111111110110111101111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111111101110111111111101111111111110110111101111111011111111111111111111111111111111101111011111100011111111110100111101111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000111111101111111111111101111111111110110011100111111011111111111111111111111111111111100111111111100011111111100100111101111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000011111100111111111111101111111111110011011110111111011111111111111111111111111111111110110111111000011111111100100111101111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000011111100001111111111011111111111110011001110111111011111111111111111111111111111100110001111111000011111111100101111100111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001111110100111111111011111111111110011101110111111011111111011111111111111111111111111111111110010011111111000101111110111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000111101110000000001111110110011111111011111111111111011100110111111011111111111111111111111111111111111111111110000011111111000001111110111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000001111101100010000001111110111100111111011111111111111111110011011111011111111111111111111111111111111111111111110000011111111000001111110111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000011111001100001000001111110111110001111111111111111111111111000011111001111111111111111111111111111111111111111110100011111110000011111110111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111110011111100110111111111111111111111110011111000111111111111111111111111111111111111111110000011111110001011111110111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000011100001000000000000111111011111110000111111111111111111111111011111000111111111111111111111111111111111111111110010011111110001011111110111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000010111111011111111100111111111111111111111111101111000111111111111111111111111111111111111111110010111111101000011111110111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000011000100000000000000111111011111111110011111111111111111111111101111000011111111111111111111111111111111111111110110111111101000111111110111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000011111011111111111000111111111111111111111101111000011111111111111111111111111111111111111110110111111001000111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111001111111111110011111111111111111111101111000001111111111111111111111111111111111111110110111111011000111111111011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001111111111111001111111111111111111110111010001111111111111111111111111111111111111100110111111011000111111111011111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111111111111100111111111111111111110111011001111111111111111110000011111111111111100110111110111000111111111011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110111111111111111111110111010000111111111111111111111001111111111111100100111110111000111111111011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111011111111111111111110111010000011111111111111111111101111111111111101101111101111000011111111011111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111111111111111011111111111111111111011010010011111111111111111111111111111111111001101111101110011011111111011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000000000111111111111111101111111111111111111011010000001111111111111111111111111111111111011101111011110011011111111011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110001000000000000011111111111111100001100111111111111011010000100111111111111111111111111111111110011101111011110011011111111001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110011100000000000011111111111111110000110000000000001011010000000011111111111111111111111111111110111101110111110011001111111001111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011100000000000011111111111111110000111110011111100001010000000001111111111111111111111111111101111101110111110111101111111101111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100011100000000000011111111111111110000011111001111111001000000000100111111111111111111111111111001111101101111100111101111111101111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111100000000000001111111111111111000001111110111111101100000000010001111111111111111111111110011111011001111101111100111111101111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111100000000000001111111111111111010001111111001111110100000000000000111111111111111111111000111111011011111111111110111111101111111111111111111011111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111000100000000011111111111111111001000111111100111110100000000000100001111111111111111100011111111010011111111111110111111101111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111001100000000011111111111111111101000011111110011111000000000000000000111111111111110001111111111010111111111111110111111101111111111111111111111100000011011111111111111111111111111111111110000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111001100000000011111111111111111101100011111111001111000000000000000100001111111110000111111111110001111111111111110011111110111111111111111111111111000000000000001111111111111111111111111110000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111011100000000011111111111111111111110001111111100111000000000000000000000111100000011111111111110011111111111111111011111110111111111111111111111111000000000000000000001111111111111111111111000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111011100000000001111111111111111111110001111111110011100100000000000000100000000111111111111111110011111111111111111011111110111111111111111111111111100000000000000000000000001111111111111111000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111011100000000001111111111111111111110001111111111001100000000000000000001111111111111111111111110111111111111111111011111110111111111111111111111111111000000000000000000000000001111111111110100000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000100111111100111110011100000000001111111111111111111111000111111110100100000000000000000001111111111111111111111111111111111111111111101111111011111111111111111111111111000000000000000000000000000001100000000010000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111110011100000000000000111111111111111111000111111110110010000000000000000001111111111111111111111111111111111111111111101111111011111111111111111111111111100000000000000000011111111111111111111100000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000011111101111110111100000000000000011111111111111111000111111110111010000000000000000001111111111111111111111111111111111111111111101111111011111111111111111111111111110000000000000000000001111111111111111111111100000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111001111110111100000000000000011111111111111111100111111111111110000010000000000011111111111111111111111111111111111111111111100111111011111111111111111111111111111100000000000000000000000000011111111111111111111111100000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000001111001111110111000000010000000001111111111111111100011111111111111000000000000000011111111111111111111111111111111111111111111110111111001111111111111111111111111111110000000000000000000000000000000111111111111111111111111111100000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000110011111100111000000100100000000111111111111111100011111111011111010000000000000011111111111111111111111111111111111111111111110111111101111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111100000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111100111000001000000000000011111111111111100011111111011111101000000000000011111111111111111111111111111111111111111111110111111101111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111110","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001001000000000011111111111111100011111111011111101100000000000011111111111111111111111111111111111111111111110011111101111111111111111111111111111111111111000000000000000000000000000000000000000000000000000010011111110","00000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000010000000000001111111111111100011111111011111110110000000000011111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000111111111111000001111111111111110110000100000001111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000111111111111000001111111101111110111000000000001111111111111111111111111111111111111111111111011111110111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100001000000000000000000011111111111000001111111101111111011100001000100101111111111111111111111111111111111111111111101111110111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000000100000001100000000000000000100010000000000000000001111111110000001111101111111111011100000000000000001111111111111111111111111111111111111111101111111011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000001100110000000000000000001111111110000001111101111111111001110000000000000000011111111111111111111111111111111111111101111111011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001001111000000000000000000111111100000001111101111111111101111000000000000000001111111111111111111111111111111111111100111111011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000010001111100000000000000000011111000000001111111111111111100111100000000000000000111111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000011111100000010000000000000100011111110000000000000000011110000000001111110111111111110111100000001000000000001111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000111111110011000000100000001001011111111001000000000000001100000000000111110111111111110111110000000001100000000111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000111111110000001110010000010011011111111100000000000000000000000000010111110111111111110011111000000000001100000011111111111111111111111111111111110011111101111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000001111111111100111110000100000111011111111110000000000000000000100000110111110111111111111011111000000000011100001000111111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000001110011111111111100000000000000000000000110111110111111111111011111100000000111110000110001111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111001111110111111111101110000000000000000000001110111110111111111111001111100000001111110000111110011111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110111111111101110000000000000010000011110111110111111111111101111110000011111110000111111001111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110111111111101110000000010000000000011110111110111111111111101111110000011111110000111111100111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110111111111101110000000000000000000111110111110111111111111111111111000000111110000111111110111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111101111111111101110100000000010000001111110111110111111111111110111111100000011110000111111111011111111111111111111111111100111111101111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111101111111111101110010000000000000011111110111110111111111111110111111110000000000000111111111011111111111111111111111111110111111101111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111101111111111111111011000000000000111111110111110111111111111111111111111000000000000011111111101111111111111111111111111110111111101111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111101111111111111111011000000000001111111110111110111111111111111011111111100000000000111111111101111111111111111111111111110111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111001111111111011111011100000000001111111110111110111111111111111011111111110000000000111111111101111111111111111111111111111011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111011111111111011111011111000000011111111110111111011111111111111011111111111000000000111111111101111111111111111111111111111011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111011111111111011111001111111000111111111110111111011111111111111101111111110110000000111111111111111111111111111111111111111011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111011111111111011111101111111111111111111110111111011111111111111101111111111011000000111111111110111111111111111111111111111011111111011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111011111111111011111101111111111111111111110111111011111111111111111111111111101100001111111111110111111111111111111111111111101111111011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110111111111111011111100111111111111111111110111111011111111111111111111111111100111111111111111110111111111111111111111111111101111111101111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110111111111111011111110111111111111111111110111111011111111111111111111111111110111111111111111011111111111111111111111111111101111111101111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111110111111111110011111110011111111111111111110111111011111111111111111111111111111011111111111111100111111111111111111111111111100111111110111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111110111111111110111111111011111111111111111110111110011111111111111111111111111111101111111111111110011111111111111111111111111110111111110111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111110111111111110111111111101111111111111111110111110011111111111111111111111111111110111111111111111011111111111111111111111111110111111110111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111101111111111110111111111100111111111111111111111110101111111111111111111111111111110111111111111111001111111111111111111111111110111111111011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000011000111111111111111111111111111111111111111101111111111110111111111110001111111111111111111101101111111111111111111111111111111011111111111111101111111111111111111111111110011111111011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111101111111111110111111111111000111111111111111111101101111111111111111111111111111111101111111111111110111111111111111111111111111011111111011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111101111111111110111111111111011000000001111111111011101111111111111111111111111111111101111111111111110111111111111111111111111111011111111101111111111111111111111111111111111111111111110000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111101111111111110111111111111101110011111111111111011101111111111111111111111111111111110111111111111111011111111111111111111111111011111111101111111111111111111111111111111111111111111111100000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111011111111111110111111111111101111111111111111110011101111111111111111111111111111111110111111111111111011111111111111111111111111101111111100111111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111011111111111110111111111111100111111111111111110111101111111111111111111111111111111110111111111111111101111111111111111111111111101111111110111111111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111011111111111110111111111111110111111111111111100111101111111111111111111111111111111111011111111111111101111111111111111111111111101111111110111111111111111111111111111111111111111111111111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111011111111111111111111111111110111111111111111101111110111111111111111111111111111111111011111111111111110111111111111111111111111101111111110011111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111011111111111101111111111111111011111111111111001111110111111111111111111111111111111111011111111111111110111111111111111111111111111111111111011111111111111111111111111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110111111111111101111111111111111011111111111111011111110111111111111111111111111111111111011111111111111111011111111111111111111111110111111111011111111111111111111111111111111111111111111100000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110111111111111101111111111111111001111111111110011111110111111111111111111111111111111111011111111111111111011111111111111111111111110111111111101111111111111111111011111111111111111111111110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110111111111111101111111111111111001111111111110111111110111111111111111111111111111111111011111111111111111011111111111111111111111110111111111101111111111111111111110111111111111111111111111100000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110111111111111101111111111111111101111111111101111111110111111111111111111111111111111111111111111111111111111111111111111111111111110011111111101111111111111111111100001111111111111111111111110000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110111111111111101111111111111111100111111111111111111110111111111111111111111111111111111111111111111111111101111111111111111111111111011111111110111111111111111111100000011111111111111111111111100000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101111111111111101111111111111111100111111111111111111110111111111111111111111111111111111101111111111111111101111111111111111111111111011111111110111111111111111111000100000111111111111111111111111000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111101111111111111111111111111111111100011111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111011111111110111111111111111111000000000011111111111111111111111100000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111101111111111111111111111111111111101111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111001111111111011111111111111111000000000000111111111111111111111111000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000111111111111111111111111111101111111111111101111111111111111101111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111101111111111011111111111111110000000000000001111111111111111111111110000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111101111111111111011111111111111111101111111111111111111111011111111111111111111111111111111101111111111111111101111111111111111111111111101111111111001111111111111111000000000000000111111111111111111101111100000000000000000000000000","00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111001111111111111011111111111111111111111111111111111111111011111111111111111111111111111111101111111111111111101111111111111111111111111101111111111101111111111111111000000000000000001111111111111111111001111000000000000000000000000","00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111011111111111111011111111111111111110111111111111111111111011111111111111111111111111111111101111111111111111101111111111111111111111111101111111111101111111111111111000000000000000000011111111111111111100011110000000000000000000000","00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111100111111111111111111111111111100000000000000000000111111111111111111000111100000000000000000000","00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111110111111111110111111111111111100000000000000000000011111111111111111100001111000000000000000000","00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111111111110111111111111111110000000000000000000000111111111111111111000011100000000000000000","00000000000000000000000000000000000000000000000000000001011111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111111111110011111111111111111000000000000000000000001111111111111111100000111100000000000000","00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111011111111111111011111111111111111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111111111111011111111111111111000000000000000000000000111111111111111110000001110000000000000","00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111011111111111111011111111111111111111011111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111110011111111111001111111111111111000000000000000000000000001111111111111111000000011100000000000","00000000000000000000000000000000000000000000000000000111111111111111111111111111111111110011111111111111011111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111011111111111001111111111111111000000000000000000000000000011111111111111111000000111000000000","00000000000000000000000000000000000000000000000000001111111111111111111111111111111111110111111111111111011111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111011111111111101011111111111111000000000000000000000000000000111111111111111000000001110000000","00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111011111111111111111111011111111111111111111111111111111111111111111111111101111111111111111111101111111111111111111111111111011111111111101111111111111111000000000000000000000000000000011111111111111110000000011100000","00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111011111111111111111111011111111111111111111111111111111111111111111111111101011111111111111111101111111111111111111111111111011111111111100111011111100010000000000000000000000000000000000111111111111111000000000111000","00000000000000000000000000000000000000000000000011111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111101111111111111111111111111111001111111111110111001111100000000000000000000000000000000000000011111111111111100000000001110","00000000000000000000000000000000000000000000000111111111111111111111111111111111111111110111111111111110111111111111111111111101111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111101111111111110111100111110000000000000000000000000000000000000000111111111111111000000000011","00000000000000000000000000000000000000000000011111111111111111111110111111111111111111110111111111111110111111111111111111111101111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111101111111111110011100001111000000000000000000000000000000000000000001111111111111110000000000","00000000000000000000000000000000000000000000111111101110110000000000011111111111111111111111111111111110111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111101111111111111011110000111100000000000000000000000000000000000000000111111111111111100000000","00000000000000000000000000000000000000000001111111101100000000000000001111111111111111111111111111111110111111111111111111111101111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111100111111111111011110000011110000000000000000000000000000000000000000001111111111111110000000","00000000000000000000000000000000000000000011111111111000000000000000000101111111111111111111111111111110111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111011111111111111111111111111111110111111111111001110000001111100000000000000000000000000000000000000000011111111111111000000","00000000000000000000000000000000000000000111111000010000000000000000000001111111111111111111111111111110111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111011111111111111111111111111111110111111111111101110000000111110000000000000000000000000000000000000000001111111111111110000","00000000000000000000000000000000000000011101100000000000000000000000000001111111111111111111111111111110111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111011111111111111111111111111111110111111111111101110000000001111000000000000000000000000000000000000000000011111111111111100","00000000000000000000000000000000000000110011000000000000000000000000000001111111111111101111111111111110111111111111111111111110111111111111111111111111111111111111111111111110111111111111111111111011111111111111111111111111111110111111111111100110000000000111100000000000000000000000000000000000000000001111111111111111","00000000000000000000000000000000000011100000000000000000000000000000000001101111111111101111111111111110111111111111111111111110011111111111111111111111111111111111111111111110111111111111111111111011111111111111111111111111111110011111111111100110000000000011110000000000000000000000000000000000000000000011111111111111","00000000000000000000000000000000000110000000000000000000000000000000000001111111111111101111111111111110111111111111111111111111011111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111011111111111110100000000000001111000000000000000000000000000000000000000000000111111111111","00000000000000000000000000000000001100100000000000000000000000000000000010111111111111101111111111111110111111111111111111111111011111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111011111111111111100000000000000111100000000000000000000000000000000000000000000011111111111","00000000000000000000000000000000110000000000000000000000000000000000000111111111111111101111111111111110111111111111111111111111011111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111011111111111111110000000000000011110000000000000000000000000000000000000000000000111111111","00000000000000000000000000000000100000000000000000000000000000000000000111111111111111101111111111111110111111111111111111111111011111111111111111111111111111111111111111111101111111111111111111110111111111111111111111111111111111001111111111111111000000000000001111100000000000000000000000000000000000000000000011111111","00000000000000000000000000000010000000000000000000000000000000000000000111111111111111101111111111111110111111111111111111111111101111111111111111111111111111111111111111111001111111111111111111110111111111111111111111111111111111101111111111111111000000000000000011110000000000000000000000000000000000000000000000111111","00000000000000000000000000000000000000000000000000000000000000000000001111111111111111001111111111111110111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111110111111111111111111111111111111111101111111111111011100000000000000001111000000000000000000000000000000000000000000000001111","00000000000000000000000000000000000000000000000000000000000000000000011111111111111111011111111111111110111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111110111111111111111111111111111111111101111111111111001110000000000000000111100000000000000000000000000000000000000000000000111","00000000000000000000000000000000000000000000000000000000000000000000011111111111111111011111111111111110111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111110111111111111111111111111111111111101111111111111001111000000000000000011110000000000000000000000000000000000000000000000001","00000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111111111110111111111111111111111111110111111111111111111111111111111111111111110111111111111111111111110111111111111111111111111111111111111111111111111100111100000000000000001111000000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000001111101111111111111011111111111111110111111111111111111111111110111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100011110000000000000000111100000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000000011111011111111111111011111111111111110111111111111111111111111110111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100001111000000000000000011110000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000001111110111111111111111011111111111111110111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111100000111100000000000000001111000000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000001111101111110111111111011111111111111110111111111111111111111111111011111111111111111111111111111111111111101111111111111111111111101111111111111111111111111111111111110111111111111100000011100000000000000000111110000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000011111111111100111111100011111111111111110111111111111111111111111111011111111111111111111111111111111111111101111111111110111111111101111111111111111111111111111111111110111111111111110000001110000000000000000001111000000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000000111110011111001111111100011111111111111110111111111111111111111111111011111111111111111111111111111111111111101111111111110111111111101111111111111111111111111111111111110011111111111110000000111000000000000000000111100000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000001111110111110001111111000011111111111111110111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111110000000011100000000000000000011110000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000011111101111100001111110000011111111111111110111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111110000000001110000000000000000001111000000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000000111111011111000001111100000011111111111111110111111111111111111111111111101111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111110000000000111000000000000000000111100000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000001111110111110000001111000000011111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111110001111011111111111111000000000011100000000000000000011111000000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000011111101111100000101110000000011111111111111110111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111110000111011111111111111000000000001110000000000000000001111100000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000000111111011111000000001100000000011111111111111110111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111110000011001111111111111000000000000111000000000000000000111110000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000001111110111111000000001000000000011111111111111110111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111111111110000001001111111111111000000000000011100000000000000000011111000000000000000000000000000000000","00000000000000000000000000000000000000000000000000000011111101111110000000011000000000011111111111111110111111111111111111111111111111011111111111111111111111111111111111111111111111110111111111111111111111111111111111111111110000001001111111111111000000000000001100000000000000000001111100000000000000000000000000000000","00000000000000000100000000000000000000000000000000000111111101111100000000110000000000011111111111111110111111111111111111111111111111011111111111111111111111111111111111111111111111110111111110111111111111111111111111111111110000000001111111111111100000000000000110000000000000000000011111000000000000000000000000000000","00000000000000001000000000000000000000000000000000001111111011111000000000100000000000011111111111111110111111111111111111111111111111011111111111111111111111111111111111111111111111111111111110011111111111111101111111111111111000000001111111111111100000000000000011000000000000000000001111100000000000000000000000000000","00000000000000010000000000000000000000000000000000011111110111110000000001000000000000011111111111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111111000111111111111111000000000111111111111100000000000000001100000000000000000000111110000000000000000000000000000","00000000000000000000000000000000000000000000000000111111101111100000000010000000000000011111111111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111101000111111111111111000000000111111111111100000000000000000110000000000000000000011111000000000000000000000000000","00000000000010000000000000000000000000000000000001111111011111000000000000000000000000011111111111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111110011111111111101000011111111111111000000000111111111111100000000000000000011000000000000000000001111100000000000000000000000000","00000000000110000000000000000000000000000000000011111110111110000000000000000000000000011111111111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111011111111011111111111000000011111111111111100000000111111111111110000000000000000001100000000000000000000111110000000000000000000000000","00000000011100000000000000000000000000000000000111111101111100000000000000000000000000011111111111111110111101111111111111111111111111101111111111111111111111111111111111111111111111111011111101011111111111000000001111111111111100000000111111111111110000000000000000000110000000000000000000011111000000000000000000000000","00000000110000000000000000000000000000000000001111111001111000000000000000000000000000011111111111111110010100111111111111111111111111101111111111111111111111111111111111111111111111111011111101001111111111000000001111111111111100000000111111111111110000000000000000000111000000000000000000001111110000000000000000000000","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111","11111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101011111111111111111111111111111111111111110111111100111110111111111111111111111111111111111111111111111111111111111111111111111");
BEGIN 
	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
	   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;